-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Monday, August 01, 2016 21:44:30 W. Europe Daylight Time

